module branch_pred(
    input IF_BP_PACKET if_bp_pkt,
    input EX_BP_PACKET ex_bp_packet,
    output BP_IF_PACKET


);
