//TODO:ADD LOGIC
module stage_ex(
    input IS_EX_PACKET is_ex_reg,
    
    output EX_IC_PACKET is_packet
);
endmodule
