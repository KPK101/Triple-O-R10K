//TODO:ADD LOGIC
module stage_is(
    input RS_IS_PACKET rs_is_packet,
    input PRF_IS_PACKET prf_is_packet,
    
    output IS_PRF_PACKET is_prf_packet,
    output IS_EX_PACKET is_packet
);
endmodule
    
