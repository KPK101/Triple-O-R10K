//TODO:ADD LOGIC
module stage_ic(
    input EX_IC_PACKET ex_ic_reg,
    
    //No Need for retire packet
    output IC_ROB_PACKET ic_rob_packet
);


endmodule
